    Mac OS X            	   2   �                                           ATTR         �   _                  �   H  com.apple.macl      �     com.apple.quarantine  	$h�:I�\T�u�                                                      q/0081;649a9c33;Brave; 