    Mac OS X            	   2   }      �                                      ATTR       �   �                     �     com.apple.quarantine q/0081;649a9c33;Brave; 