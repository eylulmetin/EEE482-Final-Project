    Mac OS X            	   2  O     �                                      ATTR      �      �                       com.apple.TextEncoding          com.apple.lastuseddate#PS         H  com.apple.macl     g     com.apple.quarantine utf-8;134217984��d             	$h�:I�\T�u� 4�*V�E�≌�>#                                    q/0081;649af3bb;TextEdit; 